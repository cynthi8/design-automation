magic
tech scmos
timestamp 1
<< metal1 >>
rect 1 5 2 6
rect 1 0 2 1
<< labels >>
rlabel space 0 0 3 6 0 .
rlabel metal1 1 0 2 1 0 1
rlabel metal1 1 5 2 6 0 2
<< end >>
