magic
tech scmos
timestamp 1618006626
<< error_s >>
rect 1 6 2 8
rect 4 6 5 8
rect 8 6 9 8
rect 11 6 12 8
rect 15 6 16 8
rect 18 6 19 8
rect 22 6 23 8
rect 25 6 26 8
rect 2 5 7 6
rect 9 5 14 6
rect 16 5 21 6
rect 23 5 28 6
rect 1 1 2 3
rect 8 1 9 3
rect 11 1 12 3
rect 15 1 16 3
rect 18 1 19 3
rect 22 1 23 3
rect 25 1 26 3
rect 2 0 7 1
rect 9 0 14 1
rect 16 0 21 1
rect 23 0 28 1
rect 5 -1 7 0
rect 1 -2 2 -1
rect 4 -2 7 -1
rect 1 -4 7 -2
rect 1 -5 8 -4
rect 1 -6 5 -5
rect 7 -6 8 -5
rect 10 -6 11 -4
rect 13 -6 14 -4
rect 16 -6 17 -4
rect 2 -7 19 -6
rect 1 -11 2 -9
rect 4 -11 5 -9
rect 7 -11 8 -9
rect 10 -11 11 -9
rect 13 -11 14 -9
rect 16 -11 17 -9
rect 2 -12 19 -11
<< error_ps >>
rect 1 -17 2 -15
rect 4 -17 5 -15
rect 8 -17 9 -15
rect 11 -17 12 -15
rect 2 -18 7 -17
rect 9 -18 14 -17
rect 1 -22 2 -20
rect 4 -22 5 -20
rect 8 -22 9 -20
rect 11 -22 12 -20
rect 2 -23 7 -22
rect 9 -23 14 -22
<< metal1 >>
rect 4 -4 5 1
rect 1 -6 2 -5
<< m2contact >>
rect 1 -5 2 -4
rect 4 -5 5 -4
<< metal2 >>
rect 2 -5 4 -4
use Cell  Cell_0
timestamp 1618002388
transform 1 0 -3 0 1 -7
box 3 7 10 15
use Cell  Cell_2
timestamp 1618002388
transform -1 0 23 0 1 -7
box 3 7 10 15
use Cell  Cell_1
timestamp 1618002388
transform 1 0 4 0 -1 13
box 3 7 10 15
use Cell  Cell_3
timestamp 1618002388
transform -1 0 30 0 -1 13
box 3 7 10 15
use Cell  Cell_4
timestamp 1618002388
transform 1 0 -3 0 1 -19
box 3 7 10 15
use Feed  Feed_0
timestamp 1618002575
transform 1 0 6 0 1 -12
box 0 0 4 8
use Feed  Feed_1
timestamp 1618002575
transform 1 0 9 0 1 -12
box 0 0 4 8
use Feed  Feed_2
timestamp 1618002575
transform 1 0 12 0 1 -12
box 0 0 4 8
use Feed  Feed_3
timestamp 1618002575
transform 1 0 15 0 1 -12
box 0 0 4 8
use Cell  Cell_5
array 0 1 7 0 0 8
timestamp 1618002388
transform 1 0 -3 0 1 -30
box 3 7 10 15
<< end >>
