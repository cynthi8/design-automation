magic
tech scmos
timestamp 1
<< metal1 >>
rect 1 0 2 1
rect 4 0 5 1
rect 1 5 2 6
rect 4 5 5 6
<< labels >>
rlabel metal1 0 0 6 6 0 .
rlabel metal1 1 0 2 1 0 1
rlabel metal1 4 0 5 1 0 2
rlabel metal1 1 5 2 6 0 3
rlabel metal1 4 5 5 6 0 4
<< end >>
