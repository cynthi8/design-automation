magic
tech scmos
timestamp 1
<< metal1 >>
rect 4 8 5 11
rect 1 6 2 7
<< m2contact >>
rect 1 7 2 8
rect 4 7 5 8
<< metal2 >>
rect 2 7 4 8
use Cell  Cell_4
timestamp 1
transform 1 0 0 0 1 11
box 0 0 6 6
use Feed  Feed_0
timestamp 1
transform 1 0 6 0 1 11
box 0 0 3 6
use Feed  Feed_1
timestamp 1
transform 1 0 9 0 1 11
box 0 0 3 6
use Feed  Feed_2
timestamp 1
transform 1 0 12 0 1 11
box 0 0 3 6
use Cell  Cell_5
array 0 1 7 0 0 8
timestamp 1
transform 1 0 15 0 1 11
box 0 0 6 6
use Cell  Cell_0
timestamp 1
transform 1 0 0 0 1 0
box 0 0 6 6
use Cell  Cell_1
timestamp 1
transform 1 0 7 0 -1 6
box 0 0 6 6
use Cell  Cell_2
timestamp 1
transform -1 0 20 0 1 0
box 0 0 6 6
use Cell  Cell_3
timestamp 1
transform -1 0 27 0 -1 6
box 0 0 6 6
use Feed  Feed_3
timestamp 1
transform 1 0 27 0 1 0
box 0 0 3 6
use Cell  Cell_6
timestamp 1
transform 1 0 30 0 1 0
box 0 0 6 6
<< labels >>
flabel space 0 11 6 17 0 FreeSans 8 0 0 0 Cell4
<< end >>
